module SlowADC (
					clk,rst
					);


endmodule
